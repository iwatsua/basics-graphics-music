`include "config.svh"

module lab_top
# (
    parameter  clk_mhz       = 125,
               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height )
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

    // assign led        = '0;
       assign abcdefgh   = '0;
       assign digit      = '0;
       assign red        = '0;
       assign green      = '0;
       assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------

    // Exercise 1: Free running counter.
    // How do you change the speed of LED blinking?
    // Try different bit slices to display.

    /*localparam w_cnt = $clog2 (clk_mhz * 1000 * 10000);

    logic [w_cnt - 1:0] cnt;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            cnt <= '0;
        else
            cnt <= cnt + 1'd1;

    assign led = cnt [$left (cnt) -: w_led];*/    

    // Exercise 2: Key-controlled counter.
    // Comment out the code above.
    // Uncomment and synthesize the code below.
    // Press the key to see the counter incrementing.

    /*wire any_key = |(~key);

    logic any_key_r;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            any_key_r <= '0;
        else
            any_key_r <= any_key;

    wire any_key_pressed = ~ any_key & any_key_r;

    logic [w_led - 1:0] cnt;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            cnt <= '0;
        else if (any_key_pressed)
            cnt <= cnt + 1'd1;

    assign led = w_led' (cnt);*/


    // Change the design, for example:
    //
    // 1. One key is used to increment, another to decrement.
    wire any_key_inc = ~key[2];
    wire any_key_dec = ~key[3];    

    logic any_key_r_inc;
    logic any_key_r_dec;    

    always_ff @ (posedge clk or posedge rst)
        if (rst) begin
            any_key_r_inc <= '0;
            any_key_r_dec <= '0;
        end
        else begin
            any_key_r_inc <= any_key_inc;
            any_key_r_dec <= any_key_dec;            
        end

    wire any_key_pressed_inc = ~ any_key_inc & any_key_r_inc;
    wire any_key_pressed_dec = ~ any_key_dec & any_key_r_dec;

    logic [w_led - 1:0] cnt;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            cnt <= '0;
        else if (any_key_pressed_inc) 
            cnt <= cnt + 1'd1;
        else if (any_key_pressed_dec) 
            cnt <= cnt - 1'd1;           

    assign led = w_led' (cnt);


    // 2. Two counters controlled by different keys
    // displayed in different groups of LEDs.
    



    

endmodule
